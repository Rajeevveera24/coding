module class8(b,f);
	input [3:0]b;
	output [3:0]f;
