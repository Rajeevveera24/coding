module class2(p,a);
	input a;
	output p;
	not (b,a);
	not (p,b);
endmodule
